module com;
initial begin

end
endmodule
