module com;
initial begin
  $display("computer");
end
endmodule
